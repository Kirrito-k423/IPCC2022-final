* layer: M1,vdd net: 1
* layer: M2,vdd net: 2
* layer: M3,vdd net: 3
R0 n2_0_100000 n2_24_100000 2.110000e+00
R1 n2_24_100000 n2_48_100000 5.600000e-01
